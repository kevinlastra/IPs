

module uart_baudgen 
  #(

  )
  ( 
    // System reset and clock
    input logic rst_n,
    input logic clk,
  )


endmodule