

module tb_uart

  
  
endmodule