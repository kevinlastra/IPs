

module tb_uart
  (
    input logic rst_n,
    input logic clk
  );

  logic rx;
  logic tx;
  logic rts_n;
  logic cts_n;
  logic wakeup;
  logic rx_irq;
  logic tx_irq;

  axi4 #(.alen(32), .xlen(32), .idlen(5)) bus(.clk(clk));

  uart #(.regmap(32'h1_0000)) uart_i 
  (
    .rst_n    (rst_n),
    .clk      (clk),
    .rx       (rx),
    .tx       (tx),
    .rts_n    (rts_n),
    .cts_n    (cts_n),
    .bus      (bus),
    .wakeup   (wakeup),
    .rx_irq   (rx_irq),
    .tx_irq   (tx_irq)
  );
  
  // DEBUG 

  logic [31:0] counter;
  logic tck;
  logic reseted;

  always_comb begin
    if(reseted) begin
      bus.aw.addr = 32'h1_0000;
      bus.aw_valid = 1;
      bus.w.data = 2604;
      bus.w_valid = 1;
    end else begin
      bus.aw.addr = 32'h1_0000;
      bus.aw_valid = 0;
      bus.w.data = 2604;
      bus.w_valid = 0;
    end
  end

  always_ff @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
      reseted <= 0;
      counter <= 0;
      tck <= 0;
    end else begin
      reseted <= 1;
      counter <= counter + 1;
      if(counter >= 1302) begin
        tck <= !tck;
        counter <= 0;
      end
    end
  end

  logic [99:0] shifter, shifter_n;

  always_comb begin
    shifter_n = shifter >> 1;
    cts_n = 0;
  end

  always_ff @(posedge tck or negedge rst_n) begin
    if(!rst_n) begin
      rx <= 1;
      shifter <= {{50{1'b1}}, 12'b100010100101, {38{1'b1}}};
    end else begin
      rx <= shifter_n[0];
      shifter <= shifter_n;
    end
  end
  
endmodule
