


package cpu_parameters;

  
  localparam int xlen = 32;
  localparam int alen = 32;
  localparam int ibus_rlen = 1;

  localparam logic [alen-1:0] START_PC = 'h0001_0000;
  
endpackage
